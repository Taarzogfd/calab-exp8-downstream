module stage_2_ID (
    input  wire clk,
    input  wire reset,

    // valid / allow
    input  wire valid_1,
    output wire allow_2,
    output  reg valid_2,
    input  wire allow_3,

    input  wire valid_3,
    input  wire valid_4,
    input  wire valid_5,

    input  wire [63:0] stage_1_to_2,
    output wire        br_taken,
    output wire [31:0] br_target,

    output wire [116:0] stage_2_to_3,
    output wire [31:0]  memory_write_data,
    
    input  wire [31:0] rf_rdata1,
    input  wire [31:0] rf_rdata2,
    output wire [ 4:0] rf_raddr1,
    output wire [ 4:0] rf_raddr2,

    input  wire [ 4:0] rf_waddr_3_fwd,
    input  wire [ 4:0] rf_waddr_4_fwd,
    input  wire [ 4:0] rf_waddr_5_fwd
);

wire readygo_2;
assign readygo_2=1'b1;

assign allow_2=~exists_hazard;

//如果当前指令是分支，那么下一拍invalid
//阻塞：如果当前出现写后读冲突，那么设置invalid直到冲突消失
always @(posedge clk) begin
    if (reset) valid_2<=1'b0;
    else if (~next_valid) valid_2<=1'b0;
    else valid_2<=valid_1;
end

wire next_valid;
wire next_invalid;
assign next_invalid = br_taken && valid_2 || exists_hazard;
assign next_valid   = ~next_invalid;

reg [63:0] upstream_input;

always @(posedge clk ) begin
    if (reset) upstream_input <= 64'b0;
    if (valid_1 && allow_3)
        upstream_input <= stage_1_to_2;
end

wire [31:0] pc;
wire [31:0] inst;

assign {inst,pc}=upstream_input;

wire        br_inst;

wire [11:0] alu_op;
wire        load_op;
wire        src1_is_pc;
wire        src2_is_imm;
wire        res_from_mem;
wire        dst_is_r1;
wire        mem_we;
wire        mem_en;
wire        src_reg_is_rd;
wire [4: 0] dest;
wire [31:0] rj_value;
wire [31:0] rkd_value;
wire [31:0] imm;
wire [31:0] br_offs;
wire [31:0] jirl_offs;

wire [ 5:0] op_31_26;
wire [ 3:0] op_25_22;
wire [ 1:0] op_21_20;
wire [ 4:0] op_19_15;
wire [ 4:0] rd;
wire [ 4:0] rj;
wire [ 4:0] rk;
wire [11:0] i12;
wire [19:0] i20;
wire [15:0] i16;
wire [25:0] i26;

wire [63:0] op_31_26_d;
wire [15:0] op_25_22_d;
wire [ 3:0] op_21_20_d;
wire [31:0] op_19_15_d;

wire        inst_add_w;
wire        inst_sub_w;
wire        inst_slt;
wire        inst_sltu;
wire        inst_nor;
wire        inst_and;
wire        inst_or;
wire        inst_xor;
wire        inst_slli_w;
wire        inst_srli_w;
wire        inst_srai_w;
wire        inst_addi_w;
wire        inst_ld_w;
wire        inst_st_w;
wire        inst_jirl;
wire        inst_b;
wire        inst_bl;
wire        inst_beq;
wire        inst_bne;
wire        inst_lu12i_w;

wire        need_ui5;
wire        need_si12;
wire        need_si16;
wire        need_si20;
wire        need_si26;
wire        src2_is_4;


wire        rf_re   ; //rf read-enable
wire        rf_we   ;
wire [ 4:0] rf_waddr;
wire [31:0] rf_wdata;

// Address Forwarding 地址前递
wire fw3_addrValid; // EX阶段的指令需要写寄存器
wire fw4_addrValid; // AM阶段的指令需要写寄存器
wire fw5_addrValid; // WB阶段的指令需要写寄存器

wire fw3_raddr1_eq; // EX的 写地址 与 第1个 读地址 相同
wire fw4_raddr1_eq; // AM的 写地址 与 第1个 读地址 相同
wire fw5_raddr1_eq; // WB的 写地址 与 第1个 读地址 相同

wire fw3_raddr2_eq; // EX的 写地址 与 第2个 读地址 相同
wire fw4_raddr2_eq; // AM的 写地址 与 第2个 读地址 相同
wire fw5_raddr2_eq; // WB的 写地址 与 第2个 读地址 相同

wire fw3_hazard_1;  // 确实存在冲突
wire fw4_hazard_1;  // 确实存在冲突
wire fw5_hazard_1;  // 确实存在冲突

wire fw3_hazard_2;  // 确实存在冲突
wire fw4_hazard_2;  // 确实存在冲突
wire fw5_hazard_2;  // 确实存在冲突

wire exists_hazard;

wire [31:0] alu_src1   ;
wire [31:0] alu_src2   ;


// Instruction to opcode
assign op_31_26  = inst[31:26];
assign op_25_22  = inst[25:22];
assign op_21_20  = inst[21:20];
assign op_19_15  = inst[19:15];

// Instruction to GPR address
assign rd   = inst[ 4: 0];
assign rj   = inst[ 9: 5];
assign rk   = inst[14:10];

// Instruction to immediate number
assign i12  = inst[21:10];
assign i20  = inst[24: 5];
assign i16  = inst[25:10];
assign i26  = {inst[ 9: 0], inst[25:10]};

// 分不同的opcode段进行译码，将其翻译为独立信号
decoder_6_64 u_dec0(.in(op_31_26 ), .out(op_31_26_d ));
decoder_4_16 u_dec1(.in(op_25_22 ), .out(op_25_22_d ));
decoder_2_4  u_dec2(.in(op_21_20 ), .out(op_21_20_d ));
decoder_5_32 u_dec3(.in(op_19_15 ), .out(op_19_15_d ));


//每个指令单独翻译出一个信号，它们是one-hot的
assign inst_add_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h00];
assign inst_sub_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h02];
assign inst_slt    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h04];
assign inst_sltu   = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h05];
assign inst_nor    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h08];
assign inst_and    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h09];
assign inst_or     = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0a];
assign inst_xor    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0b];
assign inst_slli_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h01];
assign inst_srli_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h09];
assign inst_srai_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h11];
assign inst_addi_w = op_31_26_d[6'h00] & op_25_22_d[4'ha];
assign inst_ld_w   = op_31_26_d[6'h0a] & op_25_22_d[4'h2];
assign inst_st_w   = op_31_26_d[6'h0a] & op_25_22_d[4'h6];
assign inst_jirl   = op_31_26_d[6'h13];
assign inst_b      = op_31_26_d[6'h14];
assign inst_bl     = op_31_26_d[6'h15];
assign inst_beq    = op_31_26_d[6'h16];
assign inst_bne    = op_31_26_d[6'h17];
assign inst_lu12i_w= op_31_26_d[6'h05] & ~inst[25];


// 根据指令，生成aluop
assign alu_op[ 0] = inst_add_w | inst_addi_w | inst_ld_w | inst_st_w
                    | inst_jirl | inst_bl;
assign alu_op[ 1] = inst_sub_w;
assign alu_op[ 2] = inst_slt;
assign alu_op[ 3] = inst_sltu;
assign alu_op[ 4] = inst_and;
assign alu_op[ 5] = inst_nor;
assign alu_op[ 6] = inst_or;
assign alu_op[ 7] = inst_xor;
assign alu_op[ 8] = inst_slli_w;
assign alu_op[ 9] = inst_srli_w;
assign alu_op[10] = inst_srai_w;
assign alu_op[11] = inst_lu12i_w;

// 需要immediate
assign need_ui5   =  inst_slli_w | inst_srli_w | inst_srai_w;
assign need_si12  =  inst_addi_w | inst_ld_w | inst_st_w;
assign need_si16  =  inst_jirl | inst_beq | inst_bne;
assign need_si20  =  inst_lu12i_w;
assign need_si26  =  inst_b | inst_bl;
assign src2_is_4  =  inst_jirl | inst_bl;


// 数据选择：生成立即数
assign imm = src2_is_4 ? 32'h4                      :
             need_si20 ? {i20[19:0], 12'b0}         :
/*need_ui5 || need_si12*/{{20{i12[11]}}, i12[11:0]} ;

//数据选择：branch相关的offset
assign br_offs = need_si26 ? {{ 4{i26[25]}}, i26[25:0], 2'b0} :
                             {{14{i16[15]}}, i16[15:0], 2'b0} ;

assign jirl_offs = {{14{i16[15]}}, i16[15:0], 2'b0};


// SRC相关的控制信号
assign src_reg_is_rd = inst_beq | inst_bne | inst_st_w;

assign src1_is_pc    = inst_jirl | inst_bl;

assign src2_is_imm   = inst_slli_w |
                       inst_srli_w |
                       inst_srai_w |
                       inst_addi_w |
                       inst_ld_w   |
                       inst_st_w   |
                       inst_lu12i_w|
                       inst_jirl   |
                       inst_bl     ;


//GPR相关的控制信号
assign res_from_mem  = inst_ld_w;
assign dst_is_r1     = inst_bl;
        // GENERAL PURPOSE REGISTER WRITE-ENABLE
assign rf_we         = ~inst_st_w & ~inst_beq & ~inst_bne & ~inst_b; //& ~inst_bl; 
assign mem_we        = inst_st_w;
assign mem_en        = (res_from_mem || mem_we);
assign dest          = dst_is_r1 ? 5'd1 : rd;
assign rf_re         = ~inst_lu12i_w & ~inst_b & ~inst_bl;

// Forwarded Addresses - Control Signals
assign fw3_addrValid = |rf_waddr_3_fwd; // 若该阶段的rf_we=0，地址输入时直接为0
assign fw3_raddr1_eq  = (rf_waddr_3_fwd == rf_raddr1);
assign fw3_raddr2_eq  = (rf_waddr_3_fwd == rf_raddr2);
assign fw3_hazard_1   = fw3_addrValid && fw3_raddr1_eq && valid_3;
assign fw3_hazard_2   = fw3_addrValid && fw3_raddr2_eq && valid_3;

assign fw4_addrValid = |rf_waddr_4_fwd; // 若该阶段的rf_we=0，地址输入时直接为0
assign fw4_raddr1_eq  = (rf_waddr_4_fwd == rf_raddr1);
assign fw4_raddr2_eq  = (rf_waddr_4_fwd == rf_raddr2);
assign fw4_hazard_1   = fw4_addrValid && fw4_raddr1_eq && valid_4;
assign fw4_hazard_2   = fw4_addrValid && fw4_raddr2_eq && valid_4;

assign fw5_addrValid = |rf_waddr_5_fwd; // 若该阶段的rf_we=0，地址输入时直接为0
assign fw5_raddr1_eq  = (rf_waddr_5_fwd == rf_raddr1);
assign fw5_raddr2_eq  = (rf_waddr_5_fwd == rf_raddr2);
assign fw5_hazard_1   = fw5_addrValid && fw5_raddr1_eq && valid_5;
assign fw5_hazard_2   = fw5_addrValid && fw5_raddr2_eq && valid_5;

assign exists_hazard = (((fw3_hazard_1 || fw4_hazard_1 || fw5_hazard_1) && (~src1_is_pc))|| 
                        ((fw3_hazard_2 || fw4_hazard_2 || fw5_hazard_2) && (~src2_is_imm)))
                       && rf_re;


// GPR
assign rf_raddr1 = rj;
assign rf_raddr2 = src_reg_is_rd ? rd :rk;
assign rj_value  = rf_rdata1;
assign rkd_value = rf_rdata2;


assign rj_eq_rd = (rj_value == rkd_value);

// BRANCH

assign br_taken = (   inst_beq  &&  rj_eq_rd
                   || inst_bne  && !rj_eq_rd
                   || inst_jirl
                   || inst_bl
                   || inst_b
                  )&& valid_2;// && ds_valid; 手动删除
assign br_inst = inst_beq || inst_bne || inst_bl || inst_b || inst_jirl;
assign br_target = (inst_beq || inst_bne || inst_bl || inst_b) ? (pc + br_offs) :
                                                   /*inst_jirl*/ (rj_value + jirl_offs);


//ALU
assign alu_src1 = src1_is_pc  ? pc[31:0] : rj_value;
assign alu_src2 = src2_is_imm ? imm : rkd_value;

assign stage_2_to_3={rf_we,dest,res_from_mem,alu_src1,alu_src2,alu_op,mem_we,mem_en,pc};
                    // 1 +  5  +  1             +32      + 32      + 12   +  1  +  1    +32
assign memory_write_data=rkd_value;

endmodule